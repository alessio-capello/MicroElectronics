* F:\CONTROLLO VERSIONE\MICROA\MicroB\Miller\Slew.sch

* Schematics Version 9.1 - Web Update 1
* Tue Apr 21 18:40:18 2020



** Analysis setup **
.tran 0ns 100m 0 0.01m
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Slew.net"
.INC "Slew.als"


.probe


.END
