* F:\CONTROLLO VERSIONE\MICRO\MicroB\Miller\Acm.sch

* Schematics Version 9.1 - Web Update 1
* Sat Apr 25 11:43:46 2020



** Analysis setup **
.ac DEC 1000 1 800Meg
.tran 0ns 0.25 0 0.1m
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Acm.net"
.INC "Acm.als"


.probe


.END
