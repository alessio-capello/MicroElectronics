* F:\CONTROLLO VERSIONE\MICRO\MicroB\MOSN_gm\MOSN_gm.sch

* Schematics Version 9.1 - Web Update 1
* Sat Apr 25 17:36:42 2020



** Analysis setup **
.DC LIN V_Vsd 0 3.3 100m 
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "F:\CONTROLLO VERSIONE\MICROA\MicroB\MOSN_gm\MOSN_gm.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "MOSN_gm.net"
.INC "MOSN_gm.als"


.probe


.END
