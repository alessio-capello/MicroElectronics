* F:\CONTROLLO VERSIONE\MICRO\MicroB\Miller\Vcm.sch

* Schematics Version 9.1 - Web Update 1
* Fri Apr 24 15:22:59 2020



** Analysis setup **
.ac DEC 1000 1 800Meg
.STEP LIN V_V51 0 2 0.2 
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Vcm.net"
.INC "Vcm.als"


.probe


.END
