* F:\CONTROLLO VERSIONE\MICROA\MicroB\Stadio_diff\diffP.sch

* Schematics Version 9.1 - Web Update 1
* Sat Apr 18 11:44:52 2020



** Analysis setup **
.tran 0ns 1 0 0.1m
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "diffP.net"
.INC "diffP.als"


.probe


.END
