* F:\CONTROLLO VERSIONE\MICRO\MicroB\MOSP_gm\MOSP_Vds.sch

* Schematics Version 9.1 - Web Update 1
* Sat Apr 25 18:25:32 2020



** Analysis setup **
.DC LIN V_Vds 0 3.3 20m 
.tran 0ns 1 0 0.1m
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "MOSP_Vds.net"
.INC "MOSP_Vds.als"


.probe


.END
