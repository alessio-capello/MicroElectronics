* F:\CONTROLLO VERSIONE\MICROA\MicroB\MOSP_gm\MOSP_Vds.sch

* Schematics Version 9.1 - Web Update 1
* Thu Apr 16 18:36:50 2020



** Analysis setup **
.tran 0ns 1 0 0.1m
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "MOSP_Vds.net"
.INC "MOSP_Vds.als"


.probe


.END
