* F:\CONTROLLO VERSIONE\MICRO\MicroB\Miller\Open_loop.sch

* Schematics Version 9.1 - Web Update 1
* Sat Apr 25 10:25:01 2020



** Analysis setup **
.ac DEC 1000 1 800Meg
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"
.LIB "C:\Users\Fra\Desktop\MicroB\MOSN_R0.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Open_loop.net"
.INC "Open_loop.als"


.probe


.END
