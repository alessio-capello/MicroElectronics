* F:\CONTROLLO VERSIONE\MICROA\MicroB\MOSN_gm\MOSN_gm.sch

* Schematics Version 9.1 - Web Update 1
* Wed Apr 15 17:11:28 2020



** Analysis setup **
.DC LIN V_Vgs 0 3.3 100m 
.OP 
.LIB "C:\Users\Fra\Desktop\MicroB\test.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "MOSN_gm.net"
.INC "MOSN_gm.als"


.probe


.END
